module testbench();
   reg [4:0] in;
   wire	     out;
   LUT5 #(.INIT(32'h76543210)) lut5inst(.I0(in[0]), .I1(in[1]), .I2(in[2]), .I3(in[3]), .O(out));
   initial begin
      $monitor("in 0x%x, out %d", in, out);
      in = 0;
      #1;
      in = 1;
      #1;
      in = 2;
      #1;
      in = 3;
      #1;
      in = 4;
      #1;
      in = 5;
      #1;
      in = 6;
      #1;
      in = 7;
      #1;
      in = 8;
      #1;
      in = 9;
      #1;
      in = 10;
      #1;
      in = 11;
      #1;
      in = 12;
      #1;
      in = 13;
      #1;
      in = 14;
      #1;
      in = 15;
      #1;
      in = 16;
      #1;
      in = 17;
      #1;
      in = 18;
      #1;
      in = 19;
      #1;
      in = 20;
      #1;
      in = 21;
      #1;
      in = 22;
      #1;
      in = 23;
      #1;
      in = 24;
      #1;
      in = 25;
      #1;
      in = 26;
      #1;
      in = 27;
      #1;
      in = 28;
      #1;
      in = 29;
      #1;
      in = 30;
      #1;
      in = 31;
   end
endmodule
