module testbench();
   reg [5:0] in;
   wire	     out;
   LUT6 #(.INIT(64'hfed_cba98_7654_3210)) lut6inst(.I0(in[0]), .I1(in[1]), .I2(in[2]), .I3(in[3]), .I4(in[4]), .I5(in[5]), .O(out));
   initial begin
      $monitor("in 0x%x, out %d", in, out);
      in = 0;
      #1;
      in = 1;
      #1;
      in = 2;
      #1;
      in = 3;
      #1;
      in = 4;
      #1;
      in = 5;
      #1;
      in = 6;
      #1;
      in = 7;
      #1;
      in = 8;
      #1;
      in = 9;
      #1;
      in = 10;
      #1;
      in = 11;
      #1;
      in = 12;
      #1;
      in = 13;
      #1;
      in = 14;
      #1;
      in = 15;
      #1;
      in = 16;
      #1;
      in = 17;
      #1;
      in = 18;
      #1;
      in = 19;
      #1;
      in = 20;
      #1;
      in = 21;
      #1;
      in = 22;
      #1;
      in = 23;
      #1;
      in = 24;
      #1;
      in = 25;
      #1;
      in = 26;
      #1;
      in = 27;
      #1;
      in = 28;
      #1;
      in = 29;
      #1;
      in = 30;
      #1;
      in = 31;
      #1;
      in = 32;
      #1;
      in = 33;
      #1;
      in = 34;
      #1;
      in = 35;
      #1;
      in = 36;
      #1;
      in = 37;
      #1;
      in = 38;
      #1;
      in = 39;
      #1;
      in = 40;
      #1;
      in = 41;
      #1;
      in = 42;
      #1;
      in = 43;
      #1;
      in = 44;
      #1;
      in = 45;
      #1;
      in = 46;
      #1;
      in = 47;
      #1;
      in = 48;
      #1;
      in = 49;
      #1;
      in = 50;
      #1;
      in = 51;
      #1;
      in = 52;
      #1;
      in = 53;
      #1;
      in = 54;
      #1;
      in = 55;
      #1;
      in = 56;
      #1;
      in = 57;
      #1;
      in = 58;
      #1;
      in = 59;
      #1;
      in = 60;
      #1;
      in = 61;
      #1;
      in = 62;
      #1;
      in = 63;
   end
endmodule
